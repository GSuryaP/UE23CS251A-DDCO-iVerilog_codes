module not2(c,a);
input a;
output c;
assign c=~a;
endmodule